module uart_sender(
	
	clk,
	rst_n,
	baud_set,
	send_en,
	tx_done,
	data,
	tx,
	uart_state

);

	input clk;//50mhz
	input rst_n;
	input [2:0] baud_set;
	input send_en;
	input [7:0] data;
	
	output reg tx_done;
	
	output reg tx;
	output reg uart_state;
	
	reg [7:0] stable_data;


	reg [12:0] clock_count;
	reg [12:0] cnt;
	
	reg [3:0] bit_cnt;
	
	initial cnt=0;
	
	
	always@(posedge clk or negedge rst_n)//稳定数据
		if(!rst_n)
			stable_data <= 0;
		else if(send_en)
			stable_data <= data;
		else
			stable_data <= stable_data;
	
	always@(*)//根据波特率得到1bit的时钟计数值clock_count，接下来需要根据计数值产生uart_clk
		if(!rst_n)
			clock_count <= 0;
		else
			case(baud_set)
				0:clock_count = 5207;//9600
				1:clock_count = 2603;//19200
				2:clock_count = 1301;//38400
				3:clock_count = 867;//57200
				4:clock_count = 433;//115200
				default:clock_count = 5207;//9600
			endcase
		

		
			
	always@(posedge clk or negedge rst_n) //计数一个bit维持的时间
		if(!rst_n) 
			cnt <= 0;
		else if(send_en) 
			if(cnt == clock_count)
				cnt <= 0;
			else 
				cnt <= cnt + 1;
		else if(!send_en)
			cnt <= 0;
			

			
	always@(posedge clk or negedge rst_n)//计算当前发送的是第几个bit
		if(!rst_n)
			bit_cnt <= 1;
		else if(send_en) 
			if(cnt == clock_count) begin
				if(bit_cnt == 10)
					bit_cnt <= 1;
				else 
					bit_cnt <= bit_cnt + 1;
			end
			else
				bit_cnt <= bit_cnt;
		else
			bit_cnt <= 1;	
		
	
	always@(posedge clk or negedge rst_n)
		if(!rst_n)
			tx <= 0;
		else begin
			case(bit_cnt)
				1:	tx = 1'b0;  //start bit
				2: tx = stable_data[0];
				3: tx = stable_data[1];
				4: tx = stable_data[2];
				5: tx = stable_data[3];
				6: tx = stable_data[4];
				7: tx = stable_data[5];
				8: tx = stable_data[6];
				9: tx = stable_data[7];
				10: tx = 1'b1; // stop bit
				default: tx = 1'b1;
			endcase
		end
		
	always@(posedge clk or negedge rst_n)
		if(!rst_n)
			tx_done <= 0;
		else if (cnt == clock_count && bit_cnt == 10)
			tx_done <= 1;
		else if (cnt == 0)
			tx_done <= 0;
			
	always@(posedge clk or negedge rst_n)
		if(!rst_n)
			uart_state <= 0;
		else if(send_en)
			uart_state <= 1;
		else if (cnt == clock_count)
			uart_state <= 0;
					
endmodule