module matrix_keyboard();



endmodule