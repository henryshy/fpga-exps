
module issp (
	source,
	probe);	

	output	[2:0]	source;
	input	[1:0]	probe;
endmodule
