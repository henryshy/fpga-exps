module uart2eeprom();


endmodule